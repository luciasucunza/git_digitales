library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity myMagCmp8 is
    Port ( a : in  STD_LOGIC_VECTOR (7 downto 0);
           b : in  STD_LOGIC_VECTOR (7 downto 0);
           igual : out  STD_LOGIC;
           aMayorB : out  STD_LOGIC;
           bMayorA : out  STD_LOGIC
			  );
end myMagCmp8;

architecture ARCH_myMagCmp8 of myMagCmp8 is

begin


end ARCH_myMagCmp8;

