library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity myDeco3_8 is
    Port ( entrada : in  STD_LOGIC_VECTOR (2 downto 0);
           salida : out  STD_LOGIC_VECTOR (7 downto 0)
			  );
end myDeco3_8;

architecture ARCH_myDeco3_8 of myDeco3_8 is

begin


end ARCH_myDeco3_8;

