library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity myEdgeCnt is
end myEdgeCnt;

architecture ARCH_myEdgeCnt of myEdgeCnt is

begin


end ARCH_myEdgeCnt;

