library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity myCoder4_2 is
    Port ( entrada : in  STD_LOGIC_VECTOR (3 downto 0);
           salida : out  STD_LOGIC_VECTOR (1 downto 0)
			  );
end myCoder4_2;

architecture ARCH_myCoder4_2 of myCoder4_2 is

begin


end ARCH_myCoder4_2;

